�� sr com.bankApp.Account.Account        L accountHolderst Ljava/lang/String;L currentBalancet Ljava/lang/Double;xr com.bankApp.People.Person        L 	firstNameq ~ L lastNameq ~ L passwordq ~ L usernameq ~ xpt Qq ~ q ~ t uniquet NO ONEsr java.lang.Double���J)k� D valuexr java.lang.Number������  xp        